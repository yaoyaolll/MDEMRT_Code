///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: test_p2s.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::ProASIC3> <Die::A3P1000> <Package::256 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module test_p2s( pdata24, pdata16, sdata24, sdata16 );

input pdata24, pdata16;
output sdata24, sdata16;

input [23:0] pdata24;
input [15:0] pdata16;

//<statements>

endmodule

